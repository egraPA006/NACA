module GPU (
    input [99:0] instr,
    input we,
    input [31:0] addr,
    input clk,
    output VGA_R,
    output VGA_B,
    output VGA_G,
    output v_sync,
    output h_sync
);
G
endmodule